module haha_1(
	input clk,
	input wire [9:0] characterPositionX,
	input wire [8:0] characterPositionY,
	input wire [9:0] drawingPositionX,
	input wire [8:0] drawingPositionY,
	output reg [2:0] rgb
);
	reg [9:0] x;
	reg [9:0] y;
	initial begin
		x = 'd0;
		y = 'd0;
	end

	always @(posedge clk) begin
		x <= (drawingPositionX - characterPositionX + 13);
		y <= (drawingPositionY - characterPositionY + 17);
		if(x==10 && y==9) begin	rgb <= 3'b100;	end
		else if(x==11 && y==9) begin	rgb <= 3'b100;	end
		else if(x==12 && y==9) begin	rgb <= 3'b100;	end
		else if(x==13 && y==9) begin	rgb <= 3'b100;	end
		else if(x==14 && y==9) begin	rgb <= 3'b100;	end
		else if(x==8 && y==10) begin	rgb <= 3'b100;	end
		else if(x==9 && y==10) begin	rgb <= 3'b100;	end
		else if(x==10 && y==10) begin	rgb <= 3'b110;	end
		else if(x==11 && y==10) begin	rgb <= 3'b111;	end
		else if(x==12 && y==10) begin	rgb <= 3'b110;	end
		else if(x==13 && y==10) begin	rgb <= 3'b110;	end
		else if(x==14 && y==10) begin	rgb <= 3'b110;	end
		else if(x==15 && y==10) begin	rgb <= 3'b110;	end
		else if(x==16 && y==10) begin	rgb <= 3'b100;	end
		else if(x==17 && y==10) begin	rgb <= 3'b100;	end
		else if(x==6 && y==11) begin	rgb <= 3'b100;	end
		else if(x==7 && y==11) begin	rgb <= 3'b110;	end
		else if(x==8 && y==11) begin	rgb <= 3'b110;	end
		else if(x==9 && y==11) begin	rgb <= 3'b110;	end
		else if(x==10 && y==11) begin	rgb <= 3'b111;	end
		else if(x==11 && y==11) begin	rgb <= 3'b111;	end
		else if(x==12 && y==11) begin	rgb <= 3'b111;	end
		else if(x==13 && y==11) begin	rgb <= 3'b111;	end
		else if(x==14 && y==11) begin	rgb <= 3'b111;	end
		else if(x==15 && y==11) begin	rgb <= 3'b111;	end
		else if(x==16 && y==11) begin	rgb <= 3'b110;	end
		else if(x==17 && y==11) begin	rgb <= 3'b110;	end
		else if(x==18 && y==11) begin	rgb <= 3'b110;	end
		else if(x==19 && y==11) begin	rgb <= 3'b100;	end
		else if(x==5 && y==12) begin	rgb <= 3'b100;	end
		else if(x==6 && y==12) begin	rgb <= 3'b110;	end
		else if(x==7 && y==12) begin	rgb <= 3'b110;	end
		else if(x==8 && y==12) begin	rgb <= 3'b110;	end
		else if(x==9 && y==12) begin	rgb <= 3'b110;	end
		else if(x==10 && y==12) begin	rgb <= 3'b110;	end
		else if(x==11 && y==12) begin	rgb <= 3'b111;	end
		else if(x==12 && y==12) begin	rgb <= 3'b111;	end
		else if(x==13 && y==12) begin	rgb <= 3'b111;	end
		else if(x==14 && y==12) begin	rgb <= 3'b110;	end
		else if(x==15 && y==12) begin	rgb <= 3'b110;	end
		else if(x==16 && y==12) begin	rgb <= 3'b110;	end
		else if(x==17 && y==12) begin	rgb <= 3'b110;	end
		else if(x==18 && y==12) begin	rgb <= 3'b110;	end
		else if(x==19 && y==12) begin	rgb <= 3'b100;	end
		else if(x==5 && y==13) begin	rgb <= 3'b100;	end
		else if(x==6 && y==13) begin	rgb <= 3'b110;	end
		else if(x==7 && y==13) begin	rgb <= 3'b110;	end
		else if(x==8 && y==13) begin	rgb <= 3'b110;	end
		else if(x==9 && y==13) begin	rgb <= 3'b110;	end
		else if(x==10 && y==13) begin	rgb <= 3'b111;	end
		else if(x==11 && y==13) begin	rgb <= 3'b111;	end
		else if(x==12 && y==13) begin	rgb <= 3'b111;	end
		else if(x==13 && y==13) begin	rgb <= 3'b111;	end
		else if(x==14 && y==13) begin	rgb <= 3'b111;	end
		else if(x==15 && y==13) begin	rgb <= 3'b110;	end
		else if(x==16 && y==13) begin	rgb <= 3'b110;	end
		else if(x==17 && y==13) begin	rgb <= 3'b110;	end
		else if(x==18 && y==13) begin	rgb <= 3'b110;	end
		else if(x==19 && y==13) begin	rgb <= 3'b100;	end
		else if(x==5 && y==14) begin	rgb <= 3'b100;	end
		else if(x==6 && y==14) begin	rgb <= 3'b100;	end
		else if(x==7 && y==14) begin	rgb <= 3'b110;	end
		else if(x==8 && y==14) begin	rgb <= 3'b110;	end
		else if(x==9 && y==14) begin	rgb <= 3'b110;	end
		else if(x==10 && y==14) begin	rgb <= 3'b111;	end
		else if(x==11 && y==14) begin	rgb <= 3'b111;	end
		else if(x==12 && y==14) begin	rgb <= 3'b111;	end
		else if(x==13 && y==14) begin	rgb <= 3'b111;	end
		else if(x==14 && y==14) begin	rgb <= 3'b111;	end
		else if(x==15 && y==14) begin	rgb <= 3'b111;	end
		else if(x==16 && y==14) begin	rgb <= 3'b110;	end
		else if(x==17 && y==14) begin	rgb <= 3'b110;	end
		else if(x==18 && y==14) begin	rgb <= 3'b110;	end
		else if(x==19 && y==14) begin	rgb <= 3'b100;	end
		else if(x==20 && y==14) begin	rgb <= 3'b100;	end
		else if(x==5 && y==15) begin	rgb <= 3'b100;	end
		else if(x==6 && y==15) begin	rgb <= 3'b100;	end
		else if(x==7 && y==15) begin	rgb <= 3'b110;	end
		else if(x==8 && y==15) begin	rgb <= 3'b110;	end
		else if(x==9 && y==15) begin	rgb <= 3'b110;	end
		else if(x==10 && y==15) begin	rgb <= 3'b111;	end
		else if(x==11 && y==15) begin	rgb <= 3'b111;	end
		else if(x==12 && y==15) begin	rgb <= 3'b111;	end
		else if(x==13 && y==15) begin	rgb <= 3'b111;	end
		else if(x==14 && y==15) begin	rgb <= 3'b111;	end
		else if(x==15 && y==15) begin	rgb <= 3'b111;	end
		else if(x==16 && y==15) begin	rgb <= 3'b110;	end
		else if(x==17 && y==15) begin	rgb <= 3'b110;	end
		else if(x==18 && y==15) begin	rgb <= 3'b110;	end
		else if(x==19 && y==15) begin	rgb <= 3'b100;	end
		else if(x==5 && y==16) begin	rgb <= 3'b100;	end
		else if(x==6 && y==16) begin	rgb <= 3'b100;	end
		else if(x==7 && y==16) begin	rgb <= 3'b100;	end
		else if(x==8 && y==16) begin	rgb <= 3'b110;	end
		else if(x==9 && y==16) begin	rgb <= 3'b110;	end
		else if(x==10 && y==16) begin	rgb <= 3'b110;	end
		else if(x==11 && y==16) begin	rgb <= 3'b111;	end
		else if(x==12 && y==16) begin	rgb <= 3'b110;	end
		else if(x==13 && y==16) begin	rgb <= 3'b111;	end
		else if(x==14 && y==16) begin	rgb <= 3'b111;	end
		else if(x==15 && y==16) begin	rgb <= 3'b110;	end
		else if(x==16 && y==16) begin	rgb <= 3'b110;	end
		else if(x==17 && y==16) begin	rgb <= 3'b110;	end
		else if(x==18 && y==16) begin	rgb <= 3'b110;	end
		else if(x==19 && y==16) begin	rgb <= 3'b100;	end
		else if(x==6 && y==17) begin	rgb <= 3'b100;	end
		else if(x==7 && y==17) begin	rgb <= 3'b100;	end
		else if(x==8 && y==17) begin	rgb <= 3'b110;	end
		else if(x==9 && y==17) begin	rgb <= 3'b110;	end
		else if(x==10 && y==17) begin	rgb <= 3'b100;	end
		else if(x==11 && y==17) begin	rgb <= 3'b100;	end
		else if(x==12 && y==17) begin	rgb <= 3'b110;	end
		else if(x==13 && y==17) begin	rgb <= 3'b100;	end
		else if(x==14 && y==17) begin	rgb <= 3'b100;	end
		else if(x==15 && y==17) begin	rgb <= 3'b111;	end
		else if(x==16 && y==17) begin	rgb <= 3'b111;	end
		else if(x==17 && y==17) begin	rgb <= 3'b100;	end
		else if(x==18 && y==17) begin	rgb <= 3'b100;	end
		else if(x==19 && y==17) begin	rgb <= 3'b100;	end
		else if(x==6 && y==18) begin	rgb <= 3'b100;	end
		else if(x==7 && y==18) begin	rgb <= 3'b100;	end
		else if(x==8 && y==18) begin	rgb <= 3'b100;	end
		else if(x==10 && y==18) begin	rgb <= 3'b100;	end
		else if(x==14 && y==18) begin	rgb <= 3'b100;	end
		else if(x==15 && y==18) begin	rgb <= 3'b100;	end
		else if(x==16 && y==18) begin	rgb <= 3'b100;	end
		else if(x==17 && y==18) begin	rgb <= 3'b100;	end
		else if(x==18 && y==18) begin	rgb <= 3'b100;	end
		else if(x==19 && y==18) begin	rgb <= 3'b100;	end
		else if(x==2 && y==19) begin	rgb <= 3'b101;	end
		else if(x==6 && y==19) begin	rgb <= 3'b100;	end
		else if(x==7 && y==19) begin	rgb <= 3'b100;	end
		else if(x==8 && y==19) begin	rgb <= 3'b100;	end
		else if(x==10 && y==19) begin	rgb <= 3'b100;	end
		else if(x==14 && y==19) begin	rgb <= 3'b100;	end
		else if(x==16 && y==19) begin	rgb <= 3'b100;	end
		else if(x==17 && y==19) begin	rgb <= 3'b100;	end
		else if(x==18 && y==19) begin	rgb <= 3'b110;	end
		else if(x==22 && y==19) begin	rgb <= 3'b101;	end
		else if(x==2 && y==20) begin	rgb <= 3'b111;	end
		else if(x==3 && y==20) begin	rgb <= 3'b100;	end
		else if(x==6 && y==20) begin	rgb <= 3'b110;	end
		else if(x==7 && y==20) begin	rgb <= 3'b110;	end
		else if(x==8 && y==20) begin	rgb <= 3'b110;	end
		else if(x==9 && y==20) begin	rgb <= 3'b110;	end
		else if(x==10 && y==20) begin	rgb <= 3'b100;	end
		else if(x==11 && y==20) begin	rgb <= 3'b100;	end
		else if(x==12 && y==20) begin	rgb <= 3'b110;	end
		else if(x==14 && y==20) begin	rgb <= 3'b110;	end
		else if(x==15 && y==20) begin	rgb <= 3'b110;	end
		else if(x==16 && y==20) begin	rgb <= 3'b110;	end
		else if(x==17 && y==20) begin	rgb <= 3'b110;	end
		else if(x==18 && y==20) begin	rgb <= 3'b110;	end
		else if(x==21 && y==20) begin	rgb <= 3'b100;	end
		else if(x==22 && y==20) begin	rgb <= 3'b100;	end
		else if(x==3 && y==21) begin	rgb <= 3'b100;	end
		else if(x==4 && y==21) begin	rgb <= 3'b100;	end
		else if(x==5 && y==21) begin	rgb <= 3'b100;	end
		else if(x==6 && y==21) begin	rgb <= 3'b100;	end
		else if(x==7 && y==21) begin	rgb <= 3'b110;	end
		else if(x==8 && y==21) begin	rgb <= 3'b110;	end
		else if(x==9 && y==21) begin	rgb <= 3'b100;	end
		else if(x==10 && y==21) begin	rgb <= 3'b100;	end
		else if(x==11 && y==21) begin	rgb <= 3'b110;	end
		else if(x==12 && y==21) begin	rgb <= 3'b111;	end
		else if(x==13 && y==21) begin	rgb <= 3'b100;	end
		else if(x==14 && y==21) begin	rgb <= 3'b100;	end
		else if(x==15 && y==21) begin	rgb <= 3'b111;	end
		else if(x==16 && y==21) begin	rgb <= 3'b110;	end
		else if(x==17 && y==21) begin	rgb <= 3'b111;	end
		else if(x==18 && y==21) begin	rgb <= 3'b110;	end
		else if(x==20 && y==21) begin	rgb <= 3'b100;	end
		else if(x==21 && y==21) begin	rgb <= 3'b100;	end
		else if(x==22 && y==21) begin	rgb <= 3'b111;	end
		else if(x==3 && y==22) begin	rgb <= 3'b100;	end
		else if(x==4 && y==22) begin	rgb <= 3'b100;	end
		else if(x==5 && y==22) begin	rgb <= 3'b100;	end
		else if(x==6 && y==22) begin	rgb <= 3'b100;	end
		else if(x==9 && y==22) begin	rgb <= 3'b100;	end
		else if(x==11 && y==22) begin	rgb <= 3'b100;	end
		else if(x==12 && y==22) begin	rgb <= 3'b100;	end
		else if(x==13 && y==22) begin	rgb <= 3'b100;	end
		else if(x==14 && y==22) begin	rgb <= 3'b100;	end
		else if(x==15 && y==22) begin	rgb <= 3'b100;	end
		else if(x==16 && y==22) begin	rgb <= 3'b100;	end
		else if(x==17 && y==22) begin	rgb <= 3'b100;	end
		else if(x==18 && y==22) begin	rgb <= 3'b100;	end
		else if(x==19 && y==22) begin	rgb <= 3'b100;	end
		else if(x==20 && y==22) begin	rgb <= 3'b100;	end
		else if(x==21 && y==22) begin	rgb <= 3'b100;	end
		else if(x==22 && y==22) begin	rgb <= 3'b001;	end
		else if(x==3 && y==23) begin	rgb <= 3'b100;	end
		else if(x==4 && y==23) begin	rgb <= 3'b100;	end
		else if(x==5 && y==23) begin	rgb <= 3'b100;	end
		else if(x==6 && y==23) begin	rgb <= 3'b100;	end
		else if(x==7 && y==23) begin	rgb <= 3'b100;	end
		else if(x==8 && y==23) begin	rgb <= 3'b100;	end
		else if(x==9 && y==23) begin	rgb <= 3'b110;	end
		else if(x==10 && y==23) begin	rgb <= 3'b100;	end
		else if(x==13 && y==23) begin	rgb <= 3'b100;	end
		else if(x==14 && y==23) begin	rgb <= 3'b100;	end
		else if(x==15 && y==23) begin	rgb <= 3'b100;	end
		else if(x==18 && y==23) begin	rgb <= 3'b100;	end
		else if(x==19 && y==23) begin	rgb <= 3'b100;	end
		else if(x==20 && y==23) begin	rgb <= 3'b100;	end
		else if(x==21 && y==23) begin	rgb <= 3'b110;	end
		else if(x==3 && y==24) begin	rgb <= 3'b111;	end
		else if(x==4 && y==24) begin	rgb <= 3'b100;	end
		else if(x==5 && y==24) begin	rgb <= 3'b100;	end
		else if(x==6 && y==24) begin	rgb <= 3'b100;	end
		else if(x==7 && y==24) begin	rgb <= 3'b100;	end
		else if(x==8 && y==24) begin	rgb <= 3'b100;	end
		else if(x==9 && y==24) begin	rgb <= 3'b100;	end
		else if(x==10 && y==24) begin	rgb <= 3'b110;	end
		else if(x==11 && y==24) begin	rgb <= 3'b100;	end
		else if(x==12 && y==24) begin	rgb <= 3'b100;	end
		else if(x==13 && y==24) begin	rgb <= 3'b111;	end
		else if(x==14 && y==24) begin	rgb <= 3'b110;	end
		else if(x==15 && y==24) begin	rgb <= 3'b110;	end
		else if(x==16 && y==24) begin	rgb <= 3'b100;	end
		else if(x==17 && y==24) begin	rgb <= 3'b100;	end
		else if(x==18 && y==24) begin	rgb <= 3'b100;	end
		else if(x==19 && y==24) begin	rgb <= 3'b100;	end
		else if(x==20 && y==24) begin	rgb <= 3'b100;	end
		else if(x==21 && y==24) begin	rgb <= 3'b111;	end
		else if(x==5 && y==25) begin	rgb <= 3'b100;	end
		else if(x==6 && y==25) begin	rgb <= 3'b110;	end
		else if(x==7 && y==25) begin	rgb <= 3'b110;	end
		else if(x==11 && y==25) begin	rgb <= 3'b100;	end
		else if(x==12 && y==25) begin	rgb <= 3'b110;	end
		else if(x==13 && y==25) begin	rgb <= 3'b100;	end
		else if(x==16 && y==25) begin	rgb <= 3'b110;	end
		else if(x==17 && y==25) begin	rgb <= 3'b110;	end
		else if(x==18 && y==25) begin	rgb <= 3'b110;	end
		else if(x==19 && y==25) begin	rgb <= 3'b100;	end
		else if(x==20 && y==25) begin	rgb <= 3'b100;	end
		else if(x==21 && y==25) begin	rgb <= 3'b111;	end
		else if(x==4 && y==26) begin	rgb <= 3'b100;	end
		else if(x==5 && y==26) begin	rgb <= 3'b100;	end
		else if(x==6 && y==26) begin	rgb <= 3'b100;	end
		else if(x==7 && y==26) begin	rgb <= 3'b110;	end
		else if(x==8 && y==26) begin	rgb <= 3'b100;	end
		else if(x==11 && y==26) begin	rgb <= 3'b100;	end
		else if(x==12 && y==26) begin	rgb <= 3'b100;	end
		else if(x==13 && y==26) begin	rgb <= 3'b100;	end
		else if(x==15 && y==26) begin	rgb <= 3'b100;	end
		else if(x==16 && y==26) begin	rgb <= 3'b110;	end
		else if(x==17 && y==26) begin	rgb <= 3'b110;	end
		else if(x==18 && y==26) begin	rgb <= 3'b100;	end
		else if(x==19 && y==26) begin	rgb <= 3'b100;	end
		else if(x==20 && y==26) begin	rgb <= 3'b111;	end
		else if(x==6 && y==27) begin	rgb <= 3'b100;	end
		else if(x==7 && y==27) begin	rgb <= 3'b100;	end
		else if(x==8 && y==27) begin	rgb <= 3'b110;	end
		else if(x==9 && y==27) begin	rgb <= 3'b110;	end
		else if(x==10 && y==27) begin	rgb <= 3'b100;	end
		else if(x==11 && y==27) begin	rgb <= 3'b100;	end
		else if(x==12 && y==27) begin	rgb <= 3'b100;	end
		else if(x==13 && y==27) begin	rgb <= 3'b100;	end
		else if(x==14 && y==27) begin	rgb <= 3'b110;	end
		else if(x==15 && y==27) begin	rgb <= 3'b110;	end
		else if(x==16 && y==27) begin	rgb <= 3'b100;	end
		else if(x==17 && y==27) begin	rgb <= 3'b100;	end
		else if(x==18 && y==27) begin	rgb <= 3'b100;	end
		else if(x==7 && y==28) begin	rgb <= 3'b100;	end
		else if(x==8 && y==28) begin	rgb <= 3'b110;	end
		else if(x==9 && y==28) begin	rgb <= 3'b110;	end
		else if(x==10 && y==28) begin	rgb <= 3'b110;	end
		else if(x==11 && y==28) begin	rgb <= 3'b110;	end
		else if(x==12 && y==28) begin	rgb <= 3'b100;	end
		else if(x==13 && y==28) begin	rgb <= 3'b110;	end
		else if(x==14 && y==28) begin	rgb <= 3'b110;	end
		else if(x==15 && y==28) begin	rgb <= 3'b110;	end
		else if(x==16 && y==28) begin	rgb <= 3'b100;	end
		else if(x==17 && y==28) begin	rgb <= 3'b100;	end
		else if(x==5 && y==29) begin	rgb <= 3'b111;	end
		else if(x==7 && y==29) begin	rgb <= 3'b100;	end
		else if(x==8 && y==29) begin	rgb <= 3'b100;	end
		else if(x==9 && y==29) begin	rgb <= 3'b110;	end
		else if(x==10 && y==29) begin	rgb <= 3'b110;	end
		else if(x==11 && y==29) begin	rgb <= 3'b111;	end
		else if(x==12 && y==29) begin	rgb <= 3'b111;	end
		else if(x==13 && y==29) begin	rgb <= 3'b111;	end
		else if(x==14 && y==29) begin	rgb <= 3'b110;	end
		else if(x==15 && y==29) begin	rgb <= 3'b110;	end
		else if(x==16 && y==29) begin	rgb <= 3'b100;	end
		else if(x==21 && y==29) begin	rgb <= 3'b111;	end
		else if(x==6 && y==30) begin	rgb <= 3'b110;	end
		else if(x==9 && y==30) begin	rgb <= 3'b100;	end
		else if(x==10 && y==30) begin	rgb <= 3'b100;	end
		else if(x==11 && y==30) begin	rgb <= 3'b100;	end
		else if(x==12 && y==30) begin	rgb <= 3'b100;	end
		else if(x==13 && y==30) begin	rgb <= 3'b100;	end
		else if(x==14 && y==30) begin	rgb <= 3'b100;	end
		else if(x==15 && y==30) begin	rgb <= 3'b100;	end
		else if(x==7 && y==31) begin	rgb <= 3'b111;	end
		else if(x==11 && y==31) begin	rgb <= 3'b100;	end
		else if(x==12 && y==31) begin	rgb <= 3'b100;	end
		else if(x==17 && y==31) begin	rgb <= 3'b001;	end
		else if(x==10 && y==32) begin	rgb <= 3'b100;	end
		else if(x==11 && y==32) begin	rgb <= 3'b100;	end
		else if(x==12 && y==32) begin	rgb <= 3'b100;	end
		else if(x==14 && y==32) begin	rgb <= 3'b100;	end
		else if(x==15 && y==32) begin	rgb <= 3'b111;	end
		else if(x==16 && y==32) begin	rgb <= 3'b111;	end
		else if(x==20 && y==32) begin	rgb <= 3'b111;	end
		else if(x==21 && y==32) begin	rgb <= 3'b111;	end
		else begin rgb <= 3'b000; end// Width: 25, Height: 33 From: C:/Users/guo/Pictures/Uplay/ha__.png
	end
endmodule
